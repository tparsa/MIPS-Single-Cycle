module Adder1 #(parameter N = 1)(input [