`timescale 1ns/1ns
module InstructionMem(input [15:0] address, output [15: 0] instruction, input rst);

  reg [15: 0] memory [0: 999];

 integer i;
  always @(posedge rst) begin
    for (i = 0; i < 1000; i = i + 1)
      memory[i] = 16'b0;
  end
  initial begin
    #700;
//    memory[0] = 16'b1000000010000000;
  //  memory[1] = 16'b1000011000000010;
    memory[0] = 16'b1000100000001000;
    memory[1] = 16'b0000010111110100;
    memory[2] = 16'b1000100100000010;
    memory[3] = 16'b0000010111110101;
    memory[4] = 16'b1000100100000010;
    memory[5] = 16'b0000010111110110;
    memory[6] = 16'b1000100100000010;

    memory[7] = 16'b0000010111110111;
    memory[8] = 16'b1000100100000010;
    memory[9] = 16'b0000010111111000;
    memory[10] = 16'b1000100100000010;
    memory[11] = 16'b0000010111111001;
    memory[12] = 16'b1000100100000010;
    memory[13] = 16'b0000010111111010;
    memory[14] = 16'b1000100100000010;
    memory[15] = 16'b0000010111111011;
    memory[16] = 16'b1000100100000010;
    memory[17] = 16'b0000010111111100;
    memory[18] = 16'b1000100100000010;
    memory[19] = 16'b0000010111111101;
    memory[20] = 16'b1000000001000000;
    memory[21] = 16'b1000010001000000;
    memory[22] = 16'b1000100001000000;
    memory[23] = 16'b1000100100000010;
    memory[24] = 16'b1000100000000010;
    memory[25] = 16'b1000110100000001;
    memory[26] = 16'b1000000010000001;
    memory[27] = 16'b1000010000001000;
    memory[28] = 16'b1000100000000001;
    memory[29] = 16'b1000011000000100;
    memory[30] = 16'b1000000010000010;
    memory[31] = 16'b1000010000000001;
    memory[32] = 16'b1000010000100000;
    memory[33] = 16'b0001000111111110;
    memory[34] = 16'b1100010100000101;
    memory[35] = 16'b1101010100001000;
    memory[36] = 16'b1110010100011111;
    memory[37] = 16'b1111010011001101;
    memory[38] = 16'b0010000000101010;
    memory[42] = 16'b1000111110000001;
    memory[43] = 16'b0100100111111111;
    memory[44] = 16'b0100100011111111;
    memory[255] = 16'b1000011110000011;
    memory[256] = 16'b1000011100000010;
    memory[257] = 16'b1100100100000101;
    memory[258] = 16'b1000011000010000;
  end
  assign instruction = memory[address];

endmodule